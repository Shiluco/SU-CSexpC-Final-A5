// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 Patches 1.02i SJ Lite Edition"
// CREATED		"Sat Jan 10 20:18:35 2026"

module sevenSegments(
	x3,
	x2,
	x1,
	x0,
	zero,
	one,
	two,
	three,
	four,
	five,
	six
);


input wire	x3;
input wire	x2;
input wire	x1;
input wire	x0;
output wire	zero;
output wire	one;
output wire	two;
output wire	three;
output wire	four;
output wire	five;
output wire	six;

wire	SYNTHESIZED_WIRE_88;
wire	SYNTHESIZED_WIRE_89;
wire	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_91;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_30;
wire	SYNTHESIZED_WIRE_31;
wire	SYNTHESIZED_WIRE_32;
wire	SYNTHESIZED_WIRE_33;
wire	SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_41;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_45;
wire	SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_57;
wire	SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_60;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_66;
wire	SYNTHESIZED_WIRE_67;
wire	SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_69;
wire	SYNTHESIZED_WIRE_70;
wire	SYNTHESIZED_WIRE_71;
wire	SYNTHESIZED_WIRE_72;
wire	SYNTHESIZED_WIRE_80;
wire	SYNTHESIZED_WIRE_81;
wire	SYNTHESIZED_WIRE_82;
wire	SYNTHESIZED_WIRE_83;
wire	SYNTHESIZED_WIRE_84;
wire	SYNTHESIZED_WIRE_85;




assign	SYNTHESIZED_WIRE_88 =  ~x3;

assign	SYNTHESIZED_WIRE_80 = SYNTHESIZED_WIRE_88 & x2 & SYNTHESIZED_WIRE_89;

assign	SYNTHESIZED_WIRE_14 = x1 & SYNTHESIZED_WIRE_90;

assign	SYNTHESIZED_WIRE_15 = SYNTHESIZED_WIRE_88 & x1;

assign	SYNTHESIZED_WIRE_9 = SYNTHESIZED_WIRE_91 & SYNTHESIZED_WIRE_89 & SYNTHESIZED_WIRE_90;

assign	SYNTHESIZED_WIRE_12 = x3 & SYNTHESIZED_WIRE_91 & SYNTHESIZED_WIRE_89;

assign	SYNTHESIZED_WIRE_13 = SYNTHESIZED_WIRE_9 | SYNTHESIZED_WIRE_10 | SYNTHESIZED_WIRE_11 | SYNTHESIZED_WIRE_12;

assign	zero = SYNTHESIZED_WIRE_13 | SYNTHESIZED_WIRE_14 | SYNTHESIZED_WIRE_15 | SYNTHESIZED_WIRE_16;

assign	SYNTHESIZED_WIRE_28 = SYNTHESIZED_WIRE_91 & SYNTHESIZED_WIRE_89;

assign	SYNTHESIZED_WIRE_30 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_29 = SYNTHESIZED_WIRE_88 & x1 & x0;

assign	SYNTHESIZED_WIRE_91 =  ~x2;

assign	SYNTHESIZED_WIRE_31 = SYNTHESIZED_WIRE_91 & x1 & SYNTHESIZED_WIRE_90;

assign	SYNTHESIZED_WIRE_32 = x3 & SYNTHESIZED_WIRE_89 & x0;

assign	SYNTHESIZED_WIRE_33 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_89 & SYNTHESIZED_WIRE_90;

assign	one = SYNTHESIZED_WIRE_28 | SYNTHESIZED_WIRE_29 | SYNTHESIZED_WIRE_30 | SYNTHESIZED_WIRE_31 | SYNTHESIZED_WIRE_32 | SYNTHESIZED_WIRE_33;

assign	SYNTHESIZED_WIRE_42 = SYNTHESIZED_WIRE_89 & x0;

assign	SYNTHESIZED_WIRE_40 = SYNTHESIZED_WIRE_88 & x2;

assign	SYNTHESIZED_WIRE_41 = x3 & SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_43 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_89;

assign	SYNTHESIZED_WIRE_89 =  ~x1;

assign	SYNTHESIZED_WIRE_44 = SYNTHESIZED_WIRE_88 & x0;

assign	SYNTHESIZED_WIRE_45 = SYNTHESIZED_WIRE_40 | SYNTHESIZED_WIRE_41 | SYNTHESIZED_WIRE_42;

assign	two = SYNTHESIZED_WIRE_43 | SYNTHESIZED_WIRE_44 | SYNTHESIZED_WIRE_45;

assign	SYNTHESIZED_WIRE_55 = SYNTHESIZED_WIRE_91 & SYNTHESIZED_WIRE_89 & SYNTHESIZED_WIRE_90;

assign	SYNTHESIZED_WIRE_57 = x3 & SYNTHESIZED_WIRE_91 & x0;

assign	SYNTHESIZED_WIRE_56 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_91 & x1;

assign	SYNTHESIZED_WIRE_58 = x2 & x1 & SYNTHESIZED_WIRE_90;

assign	SYNTHESIZED_WIRE_59 = x2 & SYNTHESIZED_WIRE_89 & x0;

assign	SYNTHESIZED_WIRE_90 =  ~x0;

assign	SYNTHESIZED_WIRE_60 = x3 & SYNTHESIZED_WIRE_89;

assign	three = SYNTHESIZED_WIRE_55 | SYNTHESIZED_WIRE_56 | SYNTHESIZED_WIRE_57 | SYNTHESIZED_WIRE_58 | SYNTHESIZED_WIRE_59 | SYNTHESIZED_WIRE_60;

assign	SYNTHESIZED_WIRE_65 = x1 & SYNTHESIZED_WIRE_90;

assign	SYNTHESIZED_WIRE_68 = x3 & x2;

assign	SYNTHESIZED_WIRE_66 = x3 & x1;

assign	SYNTHESIZED_WIRE_67 = SYNTHESIZED_WIRE_91 & SYNTHESIZED_WIRE_89 & SYNTHESIZED_WIRE_90;

assign	four = SYNTHESIZED_WIRE_65 | SYNTHESIZED_WIRE_66 | SYNTHESIZED_WIRE_67 | SYNTHESIZED_WIRE_68;

assign	five = SYNTHESIZED_WIRE_69 | SYNTHESIZED_WIRE_70 | SYNTHESIZED_WIRE_71 | SYNTHESIZED_WIRE_72;

assign	SYNTHESIZED_WIRE_69 = SYNTHESIZED_WIRE_89 & SYNTHESIZED_WIRE_90;

assign	SYNTHESIZED_WIRE_72 = SYNTHESIZED_WIRE_88 & x2;

assign	SYNTHESIZED_WIRE_70 = x3 & x1;

assign	SYNTHESIZED_WIRE_71 = x3 & SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_82 = x3 & SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_81 = x3 & x0;

assign	SYNTHESIZED_WIRE_83 = SYNTHESIZED_WIRE_91 & x1;

assign	SYNTHESIZED_WIRE_84 = x3 & x1;

assign	SYNTHESIZED_WIRE_85 = x1 & SYNTHESIZED_WIRE_90;

assign	six = SYNTHESIZED_WIRE_80 | SYNTHESIZED_WIRE_81 | SYNTHESIZED_WIRE_82 | SYNTHESIZED_WIRE_83 | SYNTHESIZED_WIRE_84 | SYNTHESIZED_WIRE_85;

assign	SYNTHESIZED_WIRE_10 = SYNTHESIZED_WIRE_88 & x2 & x0;

assign	SYNTHESIZED_WIRE_11 = x3 & SYNTHESIZED_WIRE_90;

assign	SYNTHESIZED_WIRE_16 = x2 & x1;


endmodule
